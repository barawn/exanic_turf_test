module xillybus_core
  (
  input  bus_clk_w,
  input  cfg_err_fatal_out_w,
  input  cfg_interrupt_msi_fail_w,
  input  cfg_interrupt_msi_sent_w,
  input [1:0] cfg_max_payload_w,
  input [2:0] cfg_max_read_req_w,
  input [3:0] cfg_rcb_status_w,
  input [63:0] m_axis_cq_tdata_w,
  input [1:0] m_axis_cq_tkeep_w,
  input  m_axis_cq_tlast_w,
  input  m_axis_cq_tvalid_w,
  input [63:0] m_axis_rc_tdata_w,
  input [1:0] m_axis_rc_tkeep_w,
  input  m_axis_rc_tlast_w,
  input  m_axis_rc_tvalid_w,
  input [5:0] pcie_rq_seq_num0_w,
  input [5:0] pcie_rq_seq_num1_w,
  input  pcie_rq_seq_num_vld0_w,
  input  pcie_rq_seq_num_vld1_w,
  input [3:0] s_axis_rq_tready_w,
  input [11:0] trn_fc_cpld_w,
  input [7:0] trn_fc_cplh_w,
  input  trn_lnk_up_n_w,
  input  trn_reset_n_w,
  input  trn_terr_drop_n_w,
  input [7:0] user_r_event_ctrl_data_w,
  input  user_r_event_ctrl_empty_w,
  input  user_r_event_ctrl_eof_w,
  input [31:0] user_r_mmresp_data_w,
  input  user_r_mmresp_empty_w,
  input  user_r_mmresp_eof_w,
  input  user_w_event_out_full_w,
  input  user_w_mmreq_full_w,
  output [3:0] GPIO_LED_w,
  output [31:0] cfg_interrupt_msi_int_w,
  output [63:0] cfg_interrupt_msi_pending_status_w,
  output  m_axis_cq_tready_w,
  output  m_axis_rc_tready_w,
  output  quiesce_w,
  output [63:0] s_axis_rq_tdata_w,
  output [1:0] s_axis_rq_tkeep_w,
  output  s_axis_rq_tlast_w,
  output [61:0] s_axis_rq_tuser_w,
  output  s_axis_rq_tvalid_w,
  output  user_r_event_ctrl_open_w,
  output  user_r_event_ctrl_rden_w,
  output  user_r_mmresp_open_w,
  output  user_r_mmresp_rden_w,
  output [31:0] user_w_event_out_data_w,
  output  user_w_event_out_open_w,
  output  user_w_event_out_wren_w,
  output [31:0] user_w_mmreq_data_w,
  output  user_w_mmreq_open_w,
  output  user_w_mmreq_wren_w
);
endmodule
